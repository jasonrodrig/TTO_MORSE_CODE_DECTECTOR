interface morse_assertions(clk , rst , dot_inp , dash_inp, char_space_inp , word_space_inp ,sout );
	
	input clk;
	input rst;
	input dot_inp;
	input dash_inp;
	input char_space_inp;
	input word_space_inp;
	input [7:0] sout; 

//assertion casses ->

endinterface
