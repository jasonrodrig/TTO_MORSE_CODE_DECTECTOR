`include "uvm_macros.svh"
package morse_pkg;
  import uvm_pkg::*;
  `include "morse_defines.sv"
  `include "morse_sequence_item.sv"
  `include "morse_sequence.sv"
  `include "morse_sequencer.sv"
  `include "morse_driver.sv"
  `include "morse_active_monitor.sv"
  `include "morse_passive_monitor.sv"
  `include "morse_active_agent.sv"
  `include "morse_passive_agent.sv"
  `include "morse_subscriber.sv"
  `include "morse_scoreboard.sv"
  `include "morse_environment.sv"
  `include "morse_test.sv"
endpackage
