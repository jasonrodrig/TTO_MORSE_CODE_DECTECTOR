`define no_of_items 5
